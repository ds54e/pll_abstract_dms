package rnm_pkg;
  timeunit 1s;
  timeprecision 1ps;

  nettype real nreal;

endpackage